b0VIM 8.0      �+{_� ;K  jerome                                  Linux                                   ~jerome/analysis/Master_LMEE/LMeeAnaFW/PlottingFW/src/jerome.h                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               utf-8U3210    #"! U                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 tpe           o                     ��������[       p              ��������J       �              ��������T                    ��������R       i             ��������Y       �             ��������Z                    ��������[       n             ��������S       �             ��������X                    ��������Z       t             ��������P       �             ��������F                    ��������L       d             ��������/       �                    4       �                    
                    ��������0                    ��������F       H             ��������9       �             ��������f       �             ��������U       -             ��������f       �             ��������f       �             ��������O       N             ��������[       �             ��������^       �             ��������i       V             ��������]       �             ��������!       	             ��������       =	             ��������       X	             ��������       t	             ��������       �	             ��������       �	             ��������       �	             ��������       �	             ��������       
             ��������        
             ��������       =
             ��������!       Y
             ��������#       z
             ��������#       �
             ��������       �
             ��������       �
             ��������       �
             ��������!                    ��������        7             ��������       W             ��������       u             ��������       �             ��������       �             ��������"       �             ��������        �             ��������                    ��������$       .             ��������       R             ��������       n             ��������"       �             ��������       �             ��������       �             ��������       �             ��������       �             ��������                    ��������       %             ��������"       9             ��������$       [             ��������                    ��������!       �             ��������       �             ��������       �             ��������       �             ��������                    ��������       .             ��������       K             ��������       h             ��������       �             ��������-       �             ��������:       �             ��������q       
             ���������       {             ���������       
             ���������       �             ��������0       $             ��������X       T             ��������e       �             ��������G                    ��������D       X             ��������i       �             ��������}                    ��������U       �             ��������R       �             ��������b       )             ��������}       �             ��������v                    ��������g       ~             ��������c       �             ��������h       H             ��������i       �                    O                                  h                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     ad     �     o       �  �  �  �  �  m  O  2    �  �  �  �  �  f  G  (  	  �  �  �  �  n  O  0    �  �  �  {  O  L     �  �  �  �  �  n  B      �
  �
  �
  b
  a
  5
  	
  
  �	  �	  �	  	  O	  #	  �  �  �  �  p  D        �  �  �  `  _  3    �  �  �  �  T  '  �  �  �  �  p  m  A      �  �  �  �  n  G  F    �  �  �  {  T  -    �  �  �  �  c  <      �  �                           "./input/LMEE_LEGO623.root",    "./input/LMEE_2017-03-16_1621.root",  //85   "./input/LMEE_2017-03-16_1041.root",   "./input/LMEE_2017-03-16_0202.root",   "./input/LMEE_2017-03-15_1701.root",    "./input/LMEE_2017-03-10_1526.root",   "./input/LMEE_2017-03-10_1245.root",  //80   "./input/LMEE_2017-03-10_0223.root",   "./input/LMEE_2017-03-09_1845.root",   "./input/LMEE_2017-03-02_1327.root",   "./input/LMEE_2017-03-01_1631.root",   "./input/LMEE_2017-03-01_0250.root",  //75   "./input/LMEE_2017-02-28_1630.root",   "./input/LMEE_2017-02-23_0202.root",    "./input/LMEE_2017-02-21_2133.root",     "./input/LMEE_2017-01-27_2230.root",   "./input/LMEE_2017-01-24_1150.root",  //70    "./input/LMEE_2017-01-16_1656.root",   "./input/LMEE_2017-01-16_1653.root",    "./input/LMEE_2017-01-13_1733.root",      "./input/LMEE_2017-01-11_1807.root", //66   "./input/LMEE_2017-01-12_0130.root", //65      "./input/LMEE_2017-01-11_0158.root", //64    "./input/LMEE_2017-01-11_0156.root", //63         "./input/LMEE_2017-01-05_0019.root", //62   "./input/LMEE_2017-01-04_1935.root", //61   "./input/LMEE_2017-01-03_1821.root", //60    "./input/LMEE_2016-12-27_1714.root", //59    "./input/LMEE_2016-12-26_0144.root", //58     "./input/LMEE_2016-12-24_0954.root", //57   "./input/LMEE_2016-12-21_0930.root", //56   "./input/LMEE_2016-12-21_0926.root", //55   "./input/LMEE_2016-12-19_1850.root", //54    "./input/LMEE_2016-12-12_1436.root", //53    "./input/LMEE_2016-12-18_1609.root", //52    "./input/LMEE_2016-12-12_0118.root", //51    "./input/LMEE_2016-12-08_1040.root", //50       "./input/LMEE_2016-12-05_0824.root", //49    "./input/LMEE_2016-12-05_0710.root", //48   "./input/LMEE_2016-12-05_0144.root", //47   "./input/LMEE_2016-12-04_2311.root", //46    "./input/LMEE_2016-11-28_1120.root", //45     "./input/LMEE_2016-11-26_0217.root", //44   "./input/LMEE_2016-11-25_1826.root", //43   "./input/LMEE_2016-11-24_1340.root", //42 ref    "./input/LMEE_2016-11-24_0136.root", //41   "./input/LMEE_2016-11-21_1306.root", //40       "./input/LMEE_2016-11-21_0035.root", //39    "./input/LMEE_2016-11-19_0254.root", //38   "./input/LMEE_2016-11-17_1602.root", //37    "./input/LMEE_2016-11-14_0150.root", //36    "./input/LMEE_2016-11-11_1359.root", //35   "./input/LMEE_2016-11-11_0226.root", //34   "./input/LMEE_2016-11-09_2338.root", //33    "./input/LMEE_2016-11-02_0212.root", //32     "./input/LMEE_2016-10-30_1109.root", //31   "./input/LMEE_2016-10-30_1106.root", //30   "./input/LMEE_2016-10-29_2244.root", //29   "./input/LMEE_2016-10-29_2239.root", //28     "./input/LMEE_2016-10-13_0159.root", //27   "./input/LMEE_2016-10-12_1633.root", //26      "./input/LMEE_2016-10-11_1253.root", //25   "./input/LMEE_2016-10-11_0207.root", //24   "./input/LMEE_2016-10-11_0203.root", //23   "./input/LMEE_23.root", //22   "./input/LMEE_22.root", //21   "./input/LMEE_21.root", //20   "./input/LMEE_20.root", //19   "./input/LMEE_19.root", //18   "./input/LMEE_18.root", //17   "./input/LMEE_17.root", //16   "./input/LMEE_16.root", //15   "./input/LMEE_15.root", //14   "./input/LMEE_14.root", //13   "./input/LMEE_13.root", //12   "./input/LMEE_12.root", //11   "./input/LMEE_11.root", //10   "./input/LMEE_10.root", //9   "./input/LMEE_9.root", //8   "./input/LMEE_8.root", //7   "./input/LMEE_7.root", //6   "./input/LMEE_6.root", //5   "./input/LMEE_5.root", //4   "./input/LMEE_4.root", //3   "./input/LMEE_3.root", //2   "./input/LMEE_2.root", //1    "./input/LMEE_1.root", //0  TString name[] = {  #include "LmBackground.h"  // input data files. make sure to edit the other strings accordingly! ad  3  [            �  �  [  Z                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     Int_t n_sconfig = sizeof(sconfig)/sizeof(*sconfig);  //SuperConfig sconfig[] = {PreFilter_0_100_18Cent,PreFilter_0_10_18Cent};//, PreFilter_0_10, PreFilter_70_100}; ad  G   �     O       �  �  �  l  K  �  �  �  �  �  �  s  4  +    �  n  ]  Z  Y  6  �  �  �  [  +        �  �  �  �    �
  �
  �
  �
  �
  �
  �
  I
  !
   
  �	  �	  	  �    �  �  �  �  U  	    �    �  C  �  �  �  5  �  �  �    0  /  �  �  �  3        �  �  �                                                                       ////SuperConfig sconfig[] = {PreFilter_0_100_1617_woPF}; //SuperConfig sconfig[] = {PreFilter_0_20};   //SuperConfig sconfig[] = {SpheroMC_0_20_all}; //  SuperConfig sconfig[] = {SpheroMC_0_20_all,SpheroMC_0_20_hard,SpheroMC_0_20_soft};  //SuperConfig sconfig[] = {Sphero_20_40_hard,Sphero_10_20_hard,Sphero_0_10_hard}; //SuperConfig sconfig[] = {Sphero_20_40_soft,Sphero_10_20_soft,Sphero_0_10_soft};  //SuperConfig sconfig[] = {Sphero_0_10_all,Sphero_0_10_hard,Sphero_0_10_soft}; //SuperConfig sconfig[] = {Sphero_0_10_hard,Sphero_0_10_soft};  //SuperConfig sconfig[] = {PreFilter_0_10_hard}; //SuperConfig sconfig[] = {PreFilter_0_10_hard,PreFilter_0_10_soft}; //  SuperConfig sconfig[] = {PreFilter_0_10_all,PreFilter_0_10_hard,PreFilter_0_10_soft}; //  SuperConfig sconfig[] = {PreFilter_0_20}; //  SuperConfig sconfig[] = {PreFilter_0_100_all}; //SuperConfig sconfig[] = {PreFilter_0_100_all, PreFilter_0_40, PreFilter_40_100}; //  SuperConfig sconfig[] = {PreFilter_0_100_all2,PreFilter_0_100_all3,PreFilter_0_100_all4}; //SuperConfig sconfig[] = {PreFilter_0_100_all, PreFilter_0_20, PreFilter_20_40, PreFilter_40_70, PreFilter_70_100}; //SuperConfig sconfig[] = {PreFilter_0_100_all, PreFilter_0_10, PreFilter_10_20, PreFilter_20_40, PreFilter_40_70, PreFilter_70_100}; //SuperConfig sconfig[] = {PreFilter_0_100_1617,PreFilter_0_100_all};//, PreFilter_0_10, PreFilter_70_100};  //  SuperConfig sconfig[] = {check_0_100_0,check_0_100_13, check_0_100_14}; //SuperConfig sconfig[] = {check_0_100_0};  //SuperConfig sconfig[] = {PreFilter_0_100_18Cent, PreFilter_0_100_18FAST, PreFilter_0_100_all};  //SuperConfig sconfig[] = {PreFilter_0_100_18Cent}; //  SuperConfig sconfig[] = {PreFilter_0_100_16f,PreFilter_0_100_17g, PreFilter_0_100_18Cent, PreFilter_0_100_18FAST}; //SuperConfig sconfig[] = {PreFilter_0_100_all,PreFilter_0_100_all3/*,PreFilter_0_100_all3*/, PreFilter_0_100_all};   SuperConfig sconfig[] = {NewPreFilter_0_100_16f,NewPreFilter_0_100_17g, NewPreFilter_0_100_18Cent, NewPreFilter_0_100_18FAST}; //SuperConfig sconfig[] = {NewPreFilter_0_100_16f,NewPreFilter_0_100_17g}; //SuperConfig sconfig[] = {NewPreFilter_0_100_18Cent, NewPreFilter_0_100_18FAST};  Double_t  kDoEtaScaling          = 1.0; Bool_t    kDoMassSlices          = kTRUE;  //kTRUE: do mass slices  kFALSE: do pair pt slices Bool_t    kUseSuperConfig        = kTRUE;    };   jpsi_list[1],4   heavyfl_files[0], heavyfl_histograms[0], 2.5,   cocktail_files[18], cocktail_files[18], cocktail_files[18], 2.155/2.13 *0.93*0.836,//.80,//1.78 0.82952 0.84   57.8, 0.99*0.95*0.99, 0.975, 1.0,   0, 20,   cconfig[64], /*mee_bins, ptee_bins,*/ LmBackground::kHybrid, SuperConfig SpheroMC_0_20_hard = {  };   jpsi_list[1],4   heavyfl_files[0], heavyfl_histograms[0], 2.5,   cocktail_files[18], cocktail_files[18], cocktail_files[18], 2.155/2.13 *0.93*1.126,//.80,//1.78 0.82952 0.84   57.8, 0.99*0.95*0.99, 0.975, 1.0,   0, 20,   cconfig[63], /*mee_bins, ptee_bins,*/ LmBackground::kHybrid, SuperConfig SpheroMC_0_20_soft = {  };   jpsi_list[1],4   heavyfl_files[0], heavyfl_histograms[0], 2.5,   cocktail_files[18], cocktail_files[18], cocktail_files[18], 2.155/2.13 *0.93,//.80,//1.78 0.82952 0.84   57.8, 0.99*0.95*0.99, 0.975, 1.0,   0, 20,   cconfig[62], /*mee_bins, ptee_bins,*/ LmBackground::kHybrid, SuperConfig SpheroMC_0_20_all = {   };   jpsi_list[1],5   heavyfl_files[0], heavyfl_histograms[0], 2.0,//1.49,   cocktail_files[17], cocktail_files[17], cocktail_files[17], 1.78/1.68*0.96,//0.9,//1.49, 0.926456 0.93   //57.8, 0.96*0.99, 0.975, 1.0,   57.8, 0.9975*0.945*0.99, 0.975, 1.0,   10, 20,   cconfig[61], /*mee_bins, ptee_bins,*/ LmBackground::kHybrid, SuperConfig SpheroMC_10_20_soft = { ad  �   �     4       �  o    �  �  D  �  �  b    �  ~  7  6  �  �  7  �
  �
  8
  �	  �	  9	  �  �  :  �  �  ,  �  �  -  �  �  �  <  �  �  �  U    �  �  \    �  �  Q  �  �  �  �  �  X  A  -                "jjung_ElectronEfficiency/pairEfficiency/reconstructedBinning/resonances/NgenPairsRecResonances:jjung_ElectronEfficiency/pairEfficiency/reconstru    "./input/efficiency/FullMC_75MeV/newGen3/Eff_CockWeighted_18c_FAST_fine_v2.root", //105   "./input/efficiency/FullMC_75MeV/newGen3/Eff_CockWeighted_18c_CENT_fine_v2.root", //104   "./input/efficiency/FullMC_75MeV/newGen3/Eff_CockWeighted_1617_fine_v2.root", //103    "./input/efficiency/FullMC_75MeV/newGen3/Eff_CockWeighted_18c_FAST_fine_v1.root", //105   "./input/efficiency/FullMC_75MeV/newGen3/Eff_CockWeighted_18c_CENT_fine_v1.root", //104   "./input/efficiency/FullMC_75MeV/newGen3/Eff_CockWeighted_1617_fine_v1.root", //103    "./input/efficiency/FullMC_75MeV/check2/Eff_CockWeighted_18_v15_2.root", //102   "./input/efficiency/FullMC_75MeV/check2/Eff_CockWeighted_18_v14_2.root", //101   "./input/efficiency/FullMC_75MeV/check2/Eff_CockWeighted_18_v13_2.root", //100   "./input/efficiency/FullMC_75MeV/check2/Eff_CockWeighted_18_v0_2.root", //99    "./input/efficiency/FullMC_75MeV/Eff_CockWeighted_17_v3.root", //98   "./input/efficiency/FullMC_75MeV/Eff_CockWeighted_16_v4.root", //97    "./input/efficiency/FullMC_75MeV/sys/Eff_CockWeighted_18cent_sys169_v6.root", //96   "./input/efficiency/FullMC_75MeV/sys/Eff_CockWeighted_18cent_sys168_v6.root", //95   "./input/efficiency/FullMC_75MeV/sys/Eff_CockWeighted_18cent_sys167_v6.root", //94   "./input/efficiency/FullMC_75MeV/sys/Eff_CockWeighted_18cent_sys166_v6.root", //93   "./input/efficiency/FullMC_75MeV/sys/Eff_CockWeighted_18cent_sys165_v6.root", //92   "./input/efficiency/FullMC_75MeV/sys/Eff_CockWeighted_18cent_sys164_v6.root", //91   "./input/efficiency/FullMC_75MeV/sys/Eff_CockWeighted_18cent_sys163_v6.root", //90  //not working   "./input/efficiency/FullMC_75MeV/sys/Eff_CockWeighted_18cent_sys162_v6.root", //89   "./input/efficiency/FullMC_75MeV/sys/Eff_CockWeighted_18cent_sys161_v6.root", //88   "./input/efficiency/FullMC_75MeV/sys/Eff_CockWeighted_18cent_sys160_v6.root", //87   "./input/efficiency/FullMC_75MeV/sys/Eff_CockWeighted_18cent_sys159_v6.root", //86   "./input/efficiency/FullMC_75MeV/sys/Eff_CockWeighted_18cent_sys158_v6.root", //85   "./input/efficiency/FullMC_75MeV/sys/Eff_CockWeighted_18cent_sys157_v6.root", //84   "./input/efficiency/FullMC_75MeV/sys/Eff_CockWeighted_18cent_sys156_v6.root", //83   "./input/efficiency/FullMC_75MeV/sys/Eff_CockWeighted_18cent_sys155_v6.root", //82   "./input/efficiency/FullMC_75MeV/sys/Eff_CockWeighted_18cent_sys154_v6.root", //81   "./input/efficiency/FullMC_75MeV/sys/Eff_CockWeighted_18cent_sys153_v6.root", //80   "./input/efficiency/FullMC_75MeV/sys/Eff_CockWeighted_18cent_sys152_v6.root", //79   "./input/efficiency/FullMC_75MeV/sys/Eff_CockWeighted_18cent_sys151_v6.root", //78   "./input/efficiency/FullMC_75MeV/sys/Eff_CockWeighted_18cent_sys150_v6.root", //77    "./input/efficiency/FullMC_75MeV/Eff_all_StatWeighted_v1.root", //76   "./input/efficiency/FullMC_75MeV/Eff_CockWeighted_18c_FAST_v6.root", //75    "./input/efficiency/FullMC_75MeV/Eff_CockWeighted_18c_CENT_v6.root", //74    "./input/efficiency/FullMC_75MeV/Eff_CockWeighted_16n17_v6.root", //73    "./input/efficiency/FullMC_75MeV/test_StatWeighted_wSDD_v1.root", //72    "./input/efficiency/FullMC_75MeV/test_StatWeighted_70-100_v5.root", //71    "./input/efficiency/FullMC_75MeV/test_StatWeighted_70-100_v2.root", //70    "./input/efficiency/FullMC_75MeV/test_StatWeighted_v7.root", //69    "./input/efficiency/FullMC_75MeV/test_2017weightedsmooth_v1.root", //68    "./input/efficiency/FullMC_75MeV/test_2018weightedsmooth_v1.root", //67    "./input/efficiency/FullMC_75MeV/test_2018weightedsmooth_fast_v1.root", //66    "./input/efficiency/FullMC_200MeV/test_2017weighted200_v2.root", //65   "./input/efficiency/FullMC_200MeV/test_2018weighted200_v2.root", //64  ad    b     
       �  �  �  �  �  �  �  �  r  b                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      "jjung_ElectronEfficiency/pairEfficiency/reconstructedBinning/resonances/NgenPairsRecResonances:jjung_ElectronEfficiency/pairEfficiency/reconstructedBinning/charm/NgenPairsRecCharm:jjung_ElectronEfficiency/pairEfficiency/reconstructedBinning/beauty/NgenPairsRecBeauty",   "NGenPairs_pt200",   "NGenPairs_pt75", TString effi_gen[] = { // name of 2D generated and reconstructed histogram };   ""   "",   "",   "", 